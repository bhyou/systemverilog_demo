/*************************************************************************
 > Copyright (C) 2021 Sangfor Ltd. All rights reserved.
 > File Name   : hello.v
 > Author      : bhyou
 > Mail        : bhyou@foxmail.com 
 > Created Time: Thu 17 Jun 2021 06:41:23 AM EDT
 ************************************************************************/
module hello;

   initial begin
      $display("\n\nhello\n");
   end
endmodule 
